//////////////////////////////////////////////////////////////////////////////////
// Company: EDA Lab, Shanghai, China
// Engineer: Hanyu Zhang
// Revision:
//          2024/11/07 created
// function:
// parameter:
//          DW: data width
// input:
// output:
// design:
// timing:
//////////////////////////////////////////////////////////////////////////////////
`ifndef __PERMUTATE_SV__
`define __PERMUTATE_SV__


`endif

